package ahb_agent_pkg;
    
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "def_file.sv"
    `include "../rtl/integration_def.sv"

    


endpackage