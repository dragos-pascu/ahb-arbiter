`timescale 1ns/1ns
package master_pkg;
    

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import integration_pkg::*;

    `include "ahb_magent_config.sv"
    `include "ahb_transaction.sv"
    `include "ahb_sequencer.sv"
    `include "ahb_master_monitor.sv"
    `include "ahb_master_driver.sv"
    `include "ahb_request.sv"
    `include "ahb_request_monitor.sv"
    `include "ahb_master_agent.sv"

    //sequences
    
    `include "sequence_lib.sv"
    


endpackage