class arbitration_coverage extends ahb_scoreboard;
    `uvm_component_utils(arbitration_coverage)

    
    

endclass
