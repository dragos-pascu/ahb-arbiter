virtual class ahb_seq extends uvm_sequence#(uvm_sequence_item);
    

    
endclass