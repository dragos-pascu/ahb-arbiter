package reset_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import integration_pkg::*;

    `include "reset_tx.sv"
    `include "reset_config.sv"
    `include "reset_sequences.sv"
    `include "reset_seqr.sv"
    `include "reset_driver.sv"
    `include "reset_agent.sv"


endpackage