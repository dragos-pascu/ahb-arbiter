/*
Signal description:

hlock : The lock signal is asserted by a master at the same time as the bus
request signal. This indicates to the arbiter that the master is
performing a number of indivisible transfers and the arbiter must
not grant any other bus master access to the bus once the first
transfer of the locked transfers has commenced. HLOCKx must
be asserted at least a cycle before the address to which it refers, in
order to prevent the arbiter from changing the grant signals.

hgrant : The grant signal is generated by the arbiter and indicates that the
appropriate master is currently the highest priority master
requesting the bus, taking into account locked transfers and
SPLIT transfers.
A master gains ownership of the address bus when HGRANTx is
HIGH and HREADY is HIGH at the rising edge of HCLK.

hmaster : The arbiter indicates which master is currently granted the bus
using the HMASTER[3:0] signals and this can be used to control
the central address and control multiplexor. The master number is
also required by SPLIT-capable slaves so that they can indicate to
the arbiter which master is able to complete a SPLIT transaction.

hmastlock : The arbiter indicates that the current transfer is part of a locked
sequence by asserting the HMASTLOCK signal, which has the
same timing as the address and control signals.

*/

import integration_pkg::*;
class ahb_transaction extends uvm_sequence_item;
        

        //transfer type
        rand transfer_t htrans;
        //address and control
        rand logic [31:0] haddr;
        rand size_t  hsize; // marimea transferului
        rand burst_t hburst; // tipul transferului
        rand rw_t hwrite; // scriere / citire
        rand logic [31:0] hwdata; // scrie data

        rand logic  hlock; // master signal
        rand logic  hbusreq; // master signal
        rand logic  hgrant; //arbiter
        rand logic[3:0] hmaster;  // arbiter
        rand logic  hsel; // decoder
        rand logic  hmastlock; // arbiter

        //slave response
        rand bit hready;
        resp_t hresp; 
        rand logic [31:0] hrdata;

    
        `uvm_object_utils_begin(ahb_transaction)
          `uvm_field_enum(transfer_t, htrans, UVM_ALL_ON)
          `uvm_field_int(haddr , UVM_ALL_ON)
          `uvm_field_enum(size_t, hsize, UVM_ALL_ON)
          `uvm_field_enum(burst_t, hburst, UVM_ALL_ON)
          `uvm_field_int(hwdata, UVM_ALL_ON)
          `uvm_field_int(hrdata, UVM_ALL_ON)
          `uvm_field_enum(rw_t,hwrite,UVM_ALL_ON)
          `uvm_field_int(hready, UVM_ALL_ON)
          `uvm_field_enum(resp_t, hresp, UVM_ALL_ON)        
        `uvm_object_utils_end

        function new(string name = "ahb_transaction");
            super.new(name);

        endfunction




endclass