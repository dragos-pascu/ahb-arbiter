class ahb_sequence_lib;
    
endclass