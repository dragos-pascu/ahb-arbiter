`timescale 1ns/1ns
package request_pkg;
    

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import integration_pkg::*;
    import ahb_seq_pkg::*;

    `include "../ahb_request_agent/ahb_request.sv"
    `include "../ahb_request_agent/config_req_agent.sv"
    `include "../ahb_request_agent/ahb_request_monitor.sv"
    `include "../ahb_request_agent/ahb_req_agent.sv"



endpackage