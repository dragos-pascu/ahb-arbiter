class ahb_env extends uvm_env;
    
    `uvm_component_utils(ahb_env)


    function new(string name="ahb_env", uvm_component parent);
        super.new(name,parent);
    endfunction

    


endclass