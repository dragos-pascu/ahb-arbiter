class ahb_slave_agent extends uvm_agent;


    


    function new(string name="ahb_slave_agent",uvm_component parent=null);
   
        super.new(name,parent);
        
    endfunction 


endclass //ahb_slave_agent extends uvm_agent