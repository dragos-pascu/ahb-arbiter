package ahb_test_pkg
    
    import uvm_pkg::*;

    `include "def_file.sv"


endpackage