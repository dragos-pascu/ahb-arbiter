class request_scoreboard extends uvm_scoreboard;
    
    `uvm_component_utils(request_scoreboard)
    `uvm_analysis_imp_decl(_predictor)
    `uvm_analysis_imp_decl(_evaluator)
    `uvm_analysis_imp_decl(_request_port)

    uvm_analysis_imp_predictor #(ahb_transaction,request_scoreboard) req_collect_predictor;
    uvm_analysis_imp_evaluator #(ahb_transaction,request_scoreboard) req_collect_evaluator;


    function new(string name = "request_scoreboard", uvm_component parent);
        super.new(name, parent);
        req_collect_predictor = new("req_collect_predictor",this);
        req_collect_evaluator =  new("req_collect_evaluator",this);
    endfunction 

    function void build_phase(uvm_phase phase);
    super.build_phase(phase);
        

    endfunction

    function void write_predictor(ahb_transaction master_item);
        
    endfunction

    function void write_evaluator(ahb_transaction slave_item);
       
    endfunction


    virtual function void check_phase(uvm_phase phase);
        

    endfunction
endclass