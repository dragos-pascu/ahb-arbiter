/*
Signal description:

hlock : The lock signal is asserted by a master at the same time as the bus
request signal. This indicates to the arbiter that the master is
performing a number of indivisible transfers and the arbiter must
not grant any other bus master access to the bus once the first
transfer of the locked transfers has commenced. HLOCKx must
be asserted at least a cycle before the haddr to which it refers, in
order to prevent the arbiter from changing the grant signals.

hgrant : The grant signal is generated by the arbiter and indicates that the
appropriate master is currently the highest priority master
requesting the bus, taking into account locked transfers and
SPLIT transfers.
A master gains ownership of the haddr bus when HGRANTx is
HIGH and HREADY is HIGH at the rising edge of HCLK.

hmaster : The arbiter indicates which master is currently granted the bus
using the HMASTER[3:0] signals and this can be used to control
the central haddr and control multiplexor. The master number is
also required by SPLIT-capable slaves so that they can indicate to
the arbiter which master is able to complete a SPLIT transaction.

hmastlock : The arbiter indicates that the current transfer is part of a locked
sequence by asserting the HMASTLOCK signal, which has the
same timing as the haddr and control signals.

*/

import integration_pkg::*;
class ahb_transaction extends uvm_sequence_item;
        

        //transfer type 
        rand transfer_t htrans[];
        //haddr and control
        rand logic [31:0] haddr[];
        rand size_t  hsize; 
        rand burst_t hburst;  
        rand rw_t hwrite; // read/write
        rand bit [31:0] hwdata[]; // 

        rand logic  hlock; // m signal to arbiter
        rand logic  hbusreq; // m signal to arbiter

        //inputs AHB master
        rand bit hready;
        resp_t hresp; 
        bit [31:0] hrdata;

        /*****Add other signals for sampling******/

    
        `uvm_object_utils_begin(ahb_transaction)
          `uvm_field_array_enum(transfer_t, htrans, UVM_ALL_ON)
          `uvm_field_array_int(haddr , UVM_ALL_ON)
          `uvm_field_enum(size_t, hsize, UVM_ALL_ON)
          `uvm_field_enum(burst_t, hburst, UVM_ALL_ON)
          `uvm_field_array_int(hwdata, UVM_ALL_ON)
          `uvm_field_int(hrdata, UVM_ALL_ON)
          `uvm_field_enum(rw_t,hwrite,UVM_ALL_ON)
          `uvm_field_int(hready, UVM_ALL_ON)
          `uvm_field_enum(resp_t, hresp, UVM_ALL_ON)
          `uvm_field_int(hlock , UVM_ALL_ON)
          `uvm_field_int(hbusreq , UVM_ALL_ON)        
        `uvm_object_utils_end

        function new(string name = "ahb_transaction");
            super.new(name);

        endfunction


        constraint address_size {
                //haddr Based on hburst and hsize
                if(hburst == SINGLE)
                        haddr.size == 1;
                if(hburst == INCR)
                        haddr.size < (1024/(2^hsize));
                if(hburst == WRAP4 || hburst == INCR4)
                        haddr.size == 4;
                if(hburst == WRAP8 || hburst == INCR8)
                        haddr.size == 8;
                if(hburst == WRAP16 || hburst == INCR16)
                        haddr.size == 16;
        }        

        constraint addr_size_limit {
                haddr.size > 0;
        }

        constraint word_boundary{
                if(hsize == HALFWORD){
                        foreach(haddr[i])
                                haddr[i][0] == 1'b0;
                }
                if(hsize == WORD){
                        foreach(haddr[i])
                                haddr[i][1:0] == 2'b0;
                }
        }

        constraint addr_val {
                if(hburst != SINGLE){
                        if(hburst == INCR || hburst == INCR4 || hburst == INCR8 || hburst == INCR16){
                                foreach(haddr[i]){
                                        if(i != 0){
                                        //ahb 2 pg 50
                                        haddr[i] == haddr[i-1] + 2**hsize;
                                        }
                                }
                        }
                }
        }          

        constraint transfer_size {
                hsize == WORD;
        }
                    
        constraint write_data {
                hwdata.size == haddr.size;
        }

        constraint nonseq_or_idle {
                if(hburst == SINGLE){
                        htrans.size == 1;
                        htrans[0] inside {IDLE, NONSEQ};
                }
        }        

        constraint burst_transfer {
                // Single transfer with no busy 
                if((haddr.size == 1) && (hburst == INCR)){
                        htrans[0] == NONSEQ; 
                }
                // Burst transfer with no busy
                else if(hburst != SINGLE){
                        htrans.size == haddr.size;
                        foreach(htrans[i]){
                                if(i == 0)
                                        htrans[i] == NONSEQ;
                                else
                                        htrans[i] == SEQ;
                        }
                } 
        }                

endclass